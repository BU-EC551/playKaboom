`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Font ROM
//////////////////////////////////////////////////////////////////////////////////
module font_rom(
	input clk,
	input [5:0] sel,		//5 bits gives up to 31 chars
	output reg [127:0] char_out
    );
	 
	always @ (posedge clk)
	begin
		char_out <= font[sel];
	end
	 
	reg [127:0] font [0:63] =  //2D array of character tiles 
		{
			
			{  8'b00000000, //0
				8'b00000000, //1
				8'b00000000, //2  
				8'b01111100, //3  *****
				8'b11000110, //4 **   **
				8'b11010110, //5 ** * **
				8'b11010110, //6 ** * **  
				8'b11010110, //7 ** * **
				8'b11010110, //8 ** * **  
				8'b11010110, //9 ** * **
				8'b11000110, //a **   **
				8'b01111100, //b  *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0
				8'b00000000, //1
				8'b00000000, //2    
				8'b00011000, //3    **
				8'b00111000, //4   ***
				8'b00011000, //5    **
				8'b00011000, //6    **
				8'b00011000, //7    **
				8'b00011000, //8    **
				8'b00011000, //9    **
				8'b00011000, //a    **
				8'b00111100, //b   ****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},

			{  8'b00000000, //0
				8'b00000000, //1
				8'b00000000, //2    
				8'b00111100, //3   ****
				8'b01100110, //4  **  **
				8'b00000010, //5       *
				8'b00000110, //6      **
				8'b00001100, //7     **
				8'b00011000, //8    **
				8'b00110000, //9   **
				8'b01100000, //a  **
				8'b01111110, //b  ******
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},		
			
			{  8'b00000000, //0
				8'b00000000, //1
				8'b00000000, //2    
				8'b00111100, //3  *****
				8'b11000110, //4 **   **
				8'b00000010, //5       *
				8'b00000110, //6      **
				8'b00001100, //7     **
				8'b00000110, //8      **
				8'b00000010, //9       *
				8'b11000110, //a **   **
				8'b00111100, //b  *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},	
		
			{  8'b00000000, //0
				8'b00000000, //1
				8'b00000000, //2    
				8'b00001110, //3     ***
				8'b00011110, //4    ****
				8'b00110110, //5   ** **
				8'b01100110, //6  **  **
				8'b11000110, //7 **   **
				8'b11111110, //8 *******
				8'b00000110, //9      **
				8'b00000110, //a      **
				8'b00000110, //b      **
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0
				8'b00000000, //1
				8'b00000000, //2    
				8'b11111110, //3 *******
				8'b11000000, //4 **   
				8'b11000000, //5 **
				8'b11000000, //6 **
				8'b11111100, //7 ******
				8'b00000110, //8      **
				8'b00000010, //9       *
				8'b11000110, //a **   **
				8'b01111100, //b  *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},	
			
			{  8'b00000000, //0
				8'b00000000, //1
				8'b00000000, //2    
				8'b01111100, //3  *****
				8'b11000110, //4 **   ** 
				8'b10000000, //5 *
				8'b10000000, //6 * 
				8'b11111100, //7 ******
				8'b11000110, //8 **   **
				8'b10000010, //9 *     *
				8'b11000110, //a **   **
				8'b01111100, //b  *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},	
			
			
			{  8'b00000000, //0
				8'b00000000, //1
				8'b00000000, //2    
				8'b11111110, //3 *******
				8'b11111110, //4 ******* 
				8'b10000010, //5       *
				8'b00000110, //6      **
				8'b00001100, //7     **
				8'b00011000, //8 	  **
				8'b00110000, //9   **
				8'b01100000, //a  **
				8'b11000000, //b ** 
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},	
			
			
			{  8'b00000000, //0
				8'b00000000, //1
				8'b00000000, //2    
				8'b01111100, //3  *****
				8'b11000110, //4 **   ** 
				8'b10000010, //5 *     *
				8'b11000110, //6 **   **
				8'b01111100, //7  *****
				8'b11000110, //8 **   **
				8'b10000010, //9 *     *
				8'b11000110, //a **   **
				8'b01111100, //b  *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},	
			
			
			{  8'b00000000, //0
				8'b00000000, //1
				8'b00000000, //2    
				8'b01111100, //3  *****
				8'b11000110, //4 **   ** 
				8'b10000010, //5 *     *
				8'b11000110, //6 **   **
				8'b01111110, //7  ******
				8'b00000010, //8       *
				8'b00000010, //9       *
				8'b11000110, //a **   **
				8'b01111100, //b  *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},	
			
			{  8'b00000000, //0	 10  6'h0A
				8'b00000000, //1
				8'b00000000, //2    
				8'b00111000, //3   ***
				8'b01101100, //4  ** **
				8'b11000110, //5 **   **
				8'b11000110, //6 **   **
				8'b11111110, //7 *******
				8'b11000110, //8 **   **
				8'b11000110, //9 **   **
				8'b11000110, //a **   **
				8'b11000110, //b **   **
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	11
				8'b00000000, //1
				8'b00000000, //2  
				8'b11111100, //3 ******
				8'b11000110, //4 **   **
				8'b11000110, //5 **   **
				8'b11000110, //6 **   **
				8'b11111110, //7 ******
				8'b11000110, //8 **   **
				8'b11000110, //9 **   **
				8'b11000110, //a **   **
				8'b11111100, //b ******
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	12
				8'b00000000, //1
				8'b00000000, //2  
				8'b01111100, //3  *****
				8'b11000110, //4 **   **
				8'b11000110, //5 **   **
				8'b11000000, //6 **     
				8'b11000000, //7 **
				8'b11000000, //8 **     
				8'b11000110, //9 **   **
				8'b11000110, //a **   **
				8'b01111100, //b  *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	13
				8'b00000000, //1
				8'b00000000, //2  
				8'b11111000, //3 *****
				8'b11001100, //4 **  **
				8'b11000110, //5 **   **
				8'b11000110, //6 **   **
				8'b11000110, //7 **   **
				8'b11000110, //8 **   **
				8'b11000110, //9 **   **
				8'b11001100, //a **  **
				8'b11111000, //b *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	14 6'h0E
				8'b00000000, //1
				8'b00000000, //2  
				8'b11111110, //3 ******
				8'b11000000, //4 **   
				8'b11000000, //5 **   
				8'b11000000, //6 **   
				8'b11111100, //7 *****
				8'b11000000, //8 **   
				8'b11000000, //9 **   
				8'b11000000, //a **   
				8'b11111100, //b ******
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	15
				8'b00000000, //1
				8'b00000000, //2  
				8'b11111110, //3 ******
				8'b11000000, //4 **   
				8'b11000000, //5 **   
				8'b11000000, //6 **   
				8'b11111100, //7 *****
				8'b11000000, //8 **   
				8'b11000000, //9 **   
				8'b11000000, //a **   
				8'b11000000, //b ** 
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	16 6'h10
				8'b00000000, //1
				8'b00000000, //2  
				8'b01111100, //3  *****
				8'b11000110, //4 **   **
				8'b11000110, //5 **   **
				8'b11000000, //6 **     
				8'b11000000, //7 **
				8'b11001110, //8 **  ***    
				8'b11000110, //9 **   **
				8'b11000110, //a **   **
				8'b01111100, //b  *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	17 6'h11
				8'b00000000, //1
				8'b00000000, //2  
				8'b11000110, //3 **   **
				8'b11000110, //4 **   **
				8'b11000110, //5 **   **
				8'b11000110, //6 **   **      
				8'b11111110, //7 *******   
				8'b11000110, //8 **   **       
				8'b11000110, //9 **   **
				8'b11000110, //a **   **
				8'b11000110, //b **   **
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	18
				8'b00000000, //1
				8'b00000000, //2  
				8'b11111110, //3 *******
				8'b00111000, //4   ***  
				8'b00111000, //5   ***  
				8'b00111000, //6   ***       
				8'b00111000, //7   ***    
				8'b00111000, //8   ***        
				8'b00111000, //9   ***  
				8'b00111000, //a   ***  
				8'b11111110, //b *******
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	19
				8'b00000000, //1
				8'b00000000, //2  
				8'b00011110, //3    ****
				8'b00001100, //4     **  
				8'b00001100, //5     **  
				8'b00001100, //6     **       
				8'b00001100, //7     **    
				8'b00001100, //8     **        
				8'b11001100, //9 **  **  
				8'b11001100, //a **  **  
				8'b01111000, //b  ****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	20
				8'b00000000, //1
				8'b00000000, //2  
				8'b11000110, //3 **   **
				8'b11000110, //4 **   **
				8'b11000110, //5 **   **
				8'b11001100, //6 **  **      
				8'b11110000, //7 ****    
				8'b11001100, //8 **  **       
				8'b11000110, //9 **   **
				8'b11000110, //a **   **
				8'b11000110, //b **   **
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	21 6'h15
				8'b00000000, //1
				8'b00000000, //2  
				8'b11000000, //3 **
				8'b11000000, //4 ** 
				8'b11000000, //5 ** 
				8'b11000000, //6 **     
				8'b11000000, //7 **   
				8'b11000000, //8 **      
				8'b11000000, //9 ** 
				8'b11111110, //a *******
				8'b11111110, //b *******
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	22 6'h16
				8'b00000000, //1
				8'b00000000, //2  
				8'b11000110, //3 **   **
				8'b11101110, //4 *** ***
				8'b11010110, //5 ** * **
				8'b11000110, //6 **   **  
				8'b11000110, //7 **   **
				8'b11000110, //8 **   **  
				8'b11000110, //9 **   **
				8'b11000110, //a **   **
				8'b11000110, //b **   **
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	23
				8'b00000000, //1
				8'b00000000, //2  
				8'b11000110, //3 **   **
				8'b11000110, //4 **   **
				8'b11100110, //5 ***  **
				8'b11110110, //6 **** **  
				8'b11011110, //7 ** ****
				8'b11001110, //8 **  ***  
				8'b11000110, //9 **   **
				8'b11000110, //a **   **
				8'b11000110, //b **   **
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	24
				8'b00000000, //1
				8'b00000000, //2  
				8'b01111100, //3  *****
				8'b11000110, //4 **   **
				8'b11000110, //5 **   **
				8'b11000110, //6 **   **  
				8'b11000110, //7 **   **
				8'b11000110, //8 **   **  
				8'b11000110, //9 **   **
				8'b11000110, //a **   **
				8'b01111100, //b  *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	25  6'h19
				8'b00000000, //1
				8'b00000000, //2  
				8'b11111100, //3 ******
				8'b11000110, //4 **   **
				8'b11000010, //5 **    *
				8'b11000110, //6 **   **
				8'b11111100, //7 ******
				8'b11000000, //8 **  
				8'b11000000, //9 **   
				8'b11000000, //a **   
				8'b11000000, //b **   
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	26 6'h1A
				8'b00000000, //1
				8'b00000000, //2  
				8'b01111100, //3  *****
				8'b11000110, //4 **   **
				8'b11000110, //5 **   **
				8'b11000110, //6 **   **  
				8'b11000110, //7 **   **
				8'b11000110, //8 **   **  
				8'b11011110, //9 ** ****
				8'b01111100, //a  *****
				8'b00000110, //b      **
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	27 6'h1B
				8'b00000000, //1
				8'b00000000, //2  
				8'b11111100, //3 ******
				8'b11000110, //4 **   **
				8'b11000010, //5 **    *
				8'b11000110, //6 **   **
				8'b11111100, //7 ******
				8'b11001100, //8 **  **
				8'b11000110, //9 **   **
				8'b11000110, //a **   **
				8'b11000110, //b **   **
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	28 6'h1C
				8'b00000000, //1
				8'b00000000, //2    
				8'b01111100, //3  *****
				8'b11000110, //4 **   ** 
				8'b10000000, //5 *     
				8'b11000000, //6 **   
				8'b01111100, //7  *****
				8'b00000110, //8      **
				8'b00000010, //9       *
				8'b11000110, //a **   **
				8'b01111100, //b  *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},	
			
			{  8'b00000000, //0	29
				8'b00000000, //1
				8'b00000000, //2  
				8'b11111110, //3 *******
				8'b00111000, //4   ***  
				8'b00111000, //5   ***  
				8'b00111000, //6   ***       
				8'b00111000, //7   ***    
				8'b00111000, //8   ***        
				8'b00111000, //9   ***  
				8'b00111000, //a   ***  
				8'b00111000, //b   ***
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	30
				8'b00000000, //1
				8'b00000000, //2  
				8'b11000110, //3 **   **
				8'b11000110, //4 **   **
				8'b11000110, //5 **   **
				8'b11000110, //6 **   **  
				8'b11000110, //7 **   **
				8'b11000110, //8 **   **  
				8'b11000110, //9 **   **
				8'b11000110, //a **   **
				8'b01111100, //b  *****
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	31
				8'b00000000, //1
				8'b00000000, //2  
				8'b11000110, //3 **   **
				8'b11000110, //4 **   **
				8'b11000110, //5 **   **
				8'b11000110, //6 **   **  
				8'b11000110, //7 **   **
				8'b11000110, //8 **   **  
				8'b01101100, //9  ** **
				8'b00111000, //a   ***
				8'b00010000, //b    * 
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	32
				8'b00000000, //1
				8'b00000000, //2  
				8'b11000110, //3 **   **
				8'b11000110, //4 **   **
				8'b11000110, //5 **   **
				8'b11000110, //6 **   **  
				8'b11000110, //7 **   **
				8'b11010110, //8 ** * **  
				8'b11010110, //9 ** * **
				8'b11101110, //a *** ***
				8'b01000100, //b  *   *  
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	33
				8'b00000000, //1
				8'b00000000, //2  
				8'b11000110, //3 **   **
				8'b11000110, //4 **   **
				8'b01101100, //5  ** **
				8'b01101100, //6  ** **  
				8'b00111000, //7   ***   
				8'b01101100, //8  ** **     
				8'b01101100, //9  ** **
				8'b11000110, //a **   **
				8'b11000110, //b **   **
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	34 6'h22
				8'b00000000, //1
				8'b00000000, //2  
				8'b11000110, //3 **   **
				8'b11000110, //4 **   **
				8'b11000110, //5 **   **
				8'b11000110, //6 **   **  
				8'b01101100, //7  ** ** 
				8'b00111000, //8   ***     
				8'b00111000, //9   *** 
				8'b00111000, //a   ***   
				8'b00111000, //b   ***  
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	35 6'h23
				8'b00000000, //1
				8'b00000000, //2  
				8'b11111110, //3 *******
				8'b11111110, //4 *******  
				8'b00000110, //5      **  
				8'b00001100, //6     **       
				8'b00011000, //7    **    
				8'b00110000, //8   **        
				8'b01100000, //9  **  
				8'b11111110, //a *******  
				8'b11111110, //b *******
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	36 6'h24
				8'b00000000, //1
				8'b00000000, //2  
				8'b00111000, //3   ***
				8'b00111000, //4   ***
				8'b00111000, //5   ***
				8'b00111000, //6   ***
				8'b00111000, //7   ***
				8'b00010000, //8    *
				8'b00000000, //9 
				8'b00111000, //a   ***
				8'b00111000, //b   ***
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	37 6'h25
				8'b00000000, //1
				8'b00000000, //2  
				8'b01111100, //3  *****
				8'b11000110, //4 **   **
				8'b11001100, //5 **   **
				8'b00011000, //6     **
				8'b00011000, //7    **
				8'b00011000, //8    **
				8'b00000000, //9    
				8'b00011000, //a    **
				8'b00011000, //b    **
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0 	38 6'h26
				8'b00000000, //1
				8'b00000000, //2  
				8'b00000000, //3   
				8'b00000000, //4   
				8'b00111000, //5   ***
				8'b00111000, //6   ***
				8'b00000000, //7   
				8'b00000000, //8    
				8'b00111000, //9   ***
				8'b00111000, //a   ***
				8'b00000000, //b   
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			},
			
			{  8'b00000000, //0	39 6'h27
				8'b00000000, //1
				8'b00000000, //2  
				8'b00000000, //3 
				8'b00000000, //4	blank
				8'b00000000, //5 
				8'b00000000, //6  
				8'b00000000, //7 
				8'b00000000, //8 
				8'b00000000, //9 
				8'b00000000, //a 
				8'b00000000, //b 
				8'b00000000, //c
				8'b00000000, //d
				8'b00000000, //e
				8'b00000000  //f
			}
			

		};
endmodule
